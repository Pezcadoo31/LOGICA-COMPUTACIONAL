
-- ABDIEL VICENCIO ANTONIO

library IEEE;
use IEEE.std_logic_1164.all;

entity MAS1_100 is 
    port ( A : in std_logic_vector (799 downto 0);
           Z : out std_logic_vector(799 downto 0));
end MAS1_100;

architecture arc of MAS1_100 is 

    component HA is
        port ( a, b : in std_logic;
               s, Cout : out std_logic
        );
    end component HA;
	 
signal C : std_logic_vector(799 downto 0);

Begin 
	
    I0 : HA port map (A(0), '1', Z(0), C(0));
    I1 : HA port map (A(1), C(0), Z(1), C(1));
    I2 : HA port map (A(2), C(1), Z(2), C(2));
    I3 : HA port map (A(3), C(2), Z(3), C(3));
    I4 : HA port map (A(4), C(3), Z(4), C(4));
    I5 : HA port map (A(5), C(4), Z(5), C(5));
    I6 : HA port map (A(6), C(5), Z(6), C(6));
    I7 : HA port map (A(7), C(6), Z(7), C(7));
    I8 : HA port map (A(8), C(7), Z(8), C(8));
    I9 : HA port map (A(9), C(8), Z(9), C(9));
	 I10 : HA port map (A(10), C(9), Z(10), C(10));
	 I11 : HA port map (A(11), C(10), Z(11), C(11));
	 I12 : HA port map (A(12), C(11), Z(12), C(12));
	 I13 : HA port map (A(13), C(12), Z(13), C(13));
	 I14 : HA port map (A(14), C(13), Z(14), C(14));
	 I15 : HA port map (A(15), C(14), Z(15), C(15));
	 I16  : HA port map (A(16), C(15), Z(16), C(16));
    I17  : HA port map (A(17), C(16), Z(17), C(17));
    I18  : HA port map (A(18), C(17), Z(18), C(18));
    I19  : HA port map (A(19), C(18), Z(19), C(19));
    I20  : HA port map (A(20), C(19), Z(20), C(20));
    I21  : HA port map (A(21), C(20), Z(21), C(21));
    I22  : HA port map (A(22), C(21), Z(22), C(22));
    I23  : HA port map (A(23), C(22), Z(23), C(23));
    I24  : HA port map (A(24), C(23), Z(24), C(24));
    I25  : HA port map (A(25), C(24), Z(25), C(25));
    I26  : HA port map (A(26), C(25), Z(26), C(26));
    I27  : HA port map (A(27), C(26), Z(27), C(27));
    I28  : HA port map (A(28), C(27), Z(28), C(28));
    I29  : HA port map (A(29), C(28), Z(29), C(29));
    I30  : HA port map (A(30), C(29), Z(30), C(30));
    I31  : HA port map (A(31), C(30), Z(31), C(31));
    I32  : HA port map (A(32), C(31), Z(32), C(32));
    I33  : HA port map (A(33), C(32), Z(33), C(33));
    I34  : HA port map (A(34), C(33), Z(34), C(34));
    I35  : HA port map (A(35), C(34), Z(35), C(35));
    I36  : HA port map (A(36), C(35), Z(36), C(36));
    I37  : HA port map (A(37), C(36), Z(37), C(37));
    I38  : HA port map (A(38), C(37), Z(38), C(38));
    I39  : HA port map (A(39), C(38), Z(39), C(39));
    I40  : HA port map (A(40), C(39), Z(40), C(40));
    I41  : HA port map (A(41), C(40), Z(41), C(41));
    I42  : HA port map (A(42), C(41), Z(42), C(42));
    I43  : HA port map (A(43), C(42), Z(43), C(43));
    I44  : HA port map (A(44), C(43), Z(44), C(44));
    I45  : HA port map (A(45), C(44), Z(45), C(45));
    I46  : HA port map (A(46), C(45), Z(46), C(46));
    I47  : HA port map (A(47), C(46), Z(47), C(47));
    I48  : HA port map (A(48), C(47), Z(48), C(48));
    I49  : HA port map (A(49), C(48), Z(49), C(49));
    I50  : HA port map (A(50), C(49), Z(50), C(50));
    I51  : HA port map (A(51), C(50), Z(51), C(51));
    I52  : HA port map (A(52), C(51), Z(52), C(52));
    I53  : HA port map (A(53), C(52), Z(53), C(53));
    I54  : HA port map (A(54), C(53), Z(54), C(54));
    I55  : HA port map (A(55), C(54), Z(55), C(55));
    I56  : HA port map (A(56), C(55), Z(56), C(56));
    I57  : HA port map (A(57), C(56), Z(57), C(57));
    I58  : HA port map (A(58), C(57), Z(58), C(58));
    I59  : HA port map (A(59), C(58), Z(59), C(59));
    I60  : HA port map (A(60), C(59), Z(60), C(60));
    I61  : HA port map (A(61), C(60), Z(61), C(61));
    I62  : HA port map (A(62), C(61), Z(62), C(62));
    I63  : HA port map (A(63), C(62), Z(63), C(63));
    I64  : HA port map (A(64), C(63), Z(64), C(64));
    I65  : HA port map (A(65), C(64), Z(65), C(65));
    I66  : HA port map (A(66), C(65), Z(66), C(66));
    I67  : HA port map (A(67), C(66), Z(67), C(67));
    I68  : HA port map (A(68), C(67), Z(68), C(68));
    I69  : HA port map (A(69), C(68), Z(69), C(69));
    I70  : HA port map (A(70), C(69), Z(70), C(70));
    I71  : HA port map (A(71), C(70), Z(71), C(71));
    I72  : HA port map (A(72), C(71), Z(72), C(72));
    I73  : HA port map (A(73), C(72), Z(73), C(73));
    I74  : HA port map (A(74), C(73), Z(74), C(74));
    I75  : HA port map (A(75), C(74), Z(75), C(75));
    I76  : HA port map (A(76), C(75), Z(76), C(76));
    I77  : HA port map (A(77), C(76), Z(77), C(77));
    I78  : HA port map (A(78), C(77), Z(78), C(78));
    I79  : HA port map (A(79), C(78), Z(79), C(79));
    I80  : HA port map (A(80), C(79), Z(80), C(80));
    I81  : HA port map (A(81), C(80), Z(81), C(81));
    I82  : HA port map (A(82), C(81), Z(82), C(82));
    I83  : HA port map (A(83), C(82), Z(83), C(83));
    I84  : HA port map (A(84), C(83), Z(84), C(84));
    I85  : HA port map (A(85), C(84), Z(85), C(85));
    I86  : HA port map (A(86), C(85), Z(86), C(86));
    I87  : HA port map (A(87), C(86), Z(87), C(87));
    I88  : HA port map (A(88), C(87), Z(88), C(88));
    I89  : HA port map (A(89), C(88), Z(89), C(89));
    I90  : HA port map (A(90), C(89), Z(90), C(90));
    I91  : HA port map (A(91), C(90), Z(91), C(91));
    I92  : HA port map (A(92), C(91), Z(92), C(92));
    I93  : HA port map (A(93), C(92), Z(93), C(93));
    I94  : HA port map (A(94), C(93), Z(94), C(94));
    I95  : HA port map (A(95), C(94), Z(95), C(95));
    I96  : HA port map (A(96), C(95), Z(96), C(96));
    I97  : HA port map (A(97), C(96), Z(97), C(97));
    I98  : HA port map (A(98), C(97), Z(98), C(98));
    I99  : HA port map (A(99), C(98), Z(99), C(99));
	 

	 I200 : HA port map (A(200), C(199), Z(200), C(200));
    I201 : HA port map (A(201), C(200), Z(201), C(201));
    I202 : HA port map (A(202), C(201), Z(202), C(202));
    I203 : HA port map (A(203), C(202), Z(203), C(203));
    I204 : HA port map (A(204), C(203), Z(204), C(204));
    I205 : HA port map (A(205), C(204), Z(205), C(205));
    I206 : HA port map (A(206), C(205), Z(206), C(206));
    I207 : HA port map (A(207), C(206), Z(207), C(207));
    I208 : HA port map (A(208), C(207), Z(208), C(208));
    I209 : HA port map (A(209), C(208), Z(209), C(209));
    I210 : HA port map (A(210), C(209), Z(210), C(210));
    I211 : HA port map (A(211), C(210), Z(211), C(211));
    I212 : HA port map (A(212), C(211), Z(212), C(212));
    I213 : HA port map (A(213), C(212), Z(213), C(213));
    I214 : HA port map (A(214), C(213), Z(214), C(214));
    I215 : HA port map (A(215), C(214), Z(215), C(215));
    I216 : HA port map (A(216), C(215), Z(216), C(216));
    I217 : HA port map (A(217), C(216), Z(217), C(217));
    I218 : HA port map (A(218), C(217), Z(218), C(218));
    I219 : HA port map (A(219), C(218), Z(219), C(219));
    I220 : HA port map (A(220), C(219), Z(220), C(220));
    I221 : HA port map (A(221), C(220), Z(221), C(221));
    I222 : HA port map (A(222), C(221), Z(222), C(222));
    I223 : HA port map (A(223), C(222), Z(223), C(223));
    I224 : HA port map (A(224), C(223), Z(224), C(224));
    I225 : HA port map (A(225), C(224), Z(225), C(225));
    I226 : HA port map (A(226), C(225), Z(226), C(226));
    I227 : HA port map (A(227), C(226), Z(227), C(227));
    I228 : HA port map (A(228), C(227), Z(228), C(228));
    I229 : HA port map (A(229), C(228), Z(229), C(229));
    I230 : HA port map (A(230), C(229), Z(230), C(230));
    I231 : HA port map (A(231), C(230), Z(231), C(231));
    I232 : HA port map (A(232), C(231), Z(232), C(232));
    I233 : HA port map (A(233), C(232), Z(233), C(233));
    I234 : HA port map (A(234), C(233), Z(234), C(234));
    I235 : HA port map (A(235), C(234), Z(235), C(235));
    I236 : HA port map (A(236), C(235), Z(236), C(236));
    I237 : HA port map (A(237), C(236), Z(237), C(237));
    I238 : HA port map (A(238), C(237), Z(238), C(238));
    I239 : HA port map (A(239), C(238), Z(239), C(239));
    I240 : HA port map (A(240), C(239), Z(240), C(240));
    I241 : HA port map (A(241), C(240), Z(241), C(241));
    I242 : HA port map (A(242), C(241), Z(242), C(242));
    I243 : HA port map (A(243), C(242), Z(243), C(243));
    I244 : HA port map (A(244), C(243), Z(244), C(244));
    I245 : HA port map (A(245), C(244), Z(245), C(245));
    I246 : HA port map (A(246), C(245), Z(246), C(246));
    I247 : HA port map (A(247), C(246), Z(247), C(247));
    I248 : HA port map (A(248), C(247), Z(248), C(248));
    I249 : HA port map (A(249), C(248), Z(249), C(249));
    I250 : HA port map (A(250), C(249), Z(250), C(250));
    I251 : HA port map (A(251), C(250), Z(251), C(251));
    I252 : HA port map (A(252), C(251), Z(252), C(252));
    I253 : HA port map (A(253), C(252), Z(253), C(253));
    I254 : HA port map (A(254), C(253), Z(254), C(254));
    I255 : HA port map (A(255), C(254), Z(255), C(255));
	 I256 : HA port map (A(256), C(255), Z(256), C(256));
    I257 : HA port map (A(257), C(256), Z(257), C(257));
	 I258 : HA port map (A(258), C(257), Z(258), C(258));
    I259 : HA port map (A(259), C(258), Z(259), C(259));
    I260 : HA port map (A(260), C(259), Z(260), C(260));
    I261 : HA port map (A(261), C(260), Z(261), C(261));
    I262 : HA port map (A(262), C(261), Z(262), C(262));
    I263 : HA port map (A(263), C(262), Z(263), C(263));
    I264 : HA port map (A(264), C(263), Z(264), C(264));
    I265 : HA port map (A(265), C(264), Z(265), C(265));
    I266 : HA port map (A(266), C(265), Z(266), C(266));
    I267 : HA port map (A(267), C(266), Z(267), C(267));
	 I268 : HA port map (A(268), C(267), Z(268), C(268));
    I269 : HA port map (A(269), C(268), Z(269), C(269));
    I270 : HA port map (A(270), C(269), Z(270), C(270));
    I271 : HA port map (A(271), C(270), Z(271), C(271));
    I272 : HA port map (A(272), C(271), Z(272), C(272));
    I273 : HA port map (A(273), C(272), Z(273), C(273));
    I274 : HA port map (A(274), C(273), Z(274), C(274));
    I275 : HA port map (A(275), C(274), Z(275), C(275));
    I276 : HA port map (A(276), C(275), Z(276), C(276));
    I277 : HA port map (A(277), C(276), Z(277), C(277));	 
	 I278 : HA port map (A(278), C(277), Z(278), C(278));
    I279 : HA port map (A(279), C(278), Z(279), C(279));
    I280 : HA port map (A(280), C(279), Z(280), C(280));
    I281 : HA port map (A(281), C(280), Z(281), C(281));
    I282 : HA port map (A(282), C(281), Z(282), C(282));
    I283 : HA port map (A(283), C(282), Z(283), C(283));
    I284 : HA port map (A(284), C(283), Z(284), C(284));
    I285 : HA port map (A(285), C(284), Z(285), C(285));
    I286 : HA port map (A(286), C(285), Z(286), C(286));
    I287 : HA port map (A(287), C(286), Z(287), C(287));
	 I288 : HA port map (A(288), C(287), Z(288), C(288));
    I289 : HA port map (A(289), C(288), Z(289), C(289));
    I290 : HA port map (A(290), C(289), Z(290), C(290));
    I291 : HA port map (A(291), C(290), Z(291), C(291));
    I292 : HA port map (A(292), C(291), Z(292), C(292));
    I293 : HA port map (A(293), C(292), Z(293), C(293));
    I294 : HA port map (A(294), C(293), Z(294), C(294));
    I295 : HA port map (A(295), C(294), Z(295), C(295));
    I296 : HA port map (A(296), C(295), Z(296), C(296));
    I297 : HA port map (A(297), C(296), Z(297), C(297));
    I298 : HA port map (A(298), C(297), Z(298), C(298));
    I299 : HA port map (A(299), C(298), Z(299), C(299));
    I300 : HA port map (A(300), C(299), Z(300), C(300));
    I301 : HA port map (A(301), C(300), Z(301), C(301));
    I302 : HA port map (A(302), C(301), Z(302), C(302));
    I303 : HA port map (A(303), C(302), Z(303), C(303));
    I304 : HA port map (A(304), C(303), Z(304), C(304));
    I305 : HA port map (A(305), C(304), Z(305), C(305));
    I306 : HA port map (A(306), C(305), Z(306), C(306));
    I307 : HA port map (A(307), C(306), Z(307), C(307)); 
	 I308 : HA port map (A(308), C(307), Z(308), C(308));
    I309 : HA port map (A(309), C(308), Z(309), C(309));
    I310 : HA port map (A(310), C(309), Z(310), C(310));
    I311 : HA port map (A(311), C(310), Z(311), C(311));
    I312 : HA port map (A(312), C(311), Z(312), C(312));
    I313 : HA port map (A(313), C(312), Z(313), C(313));
    I314 : HA port map (A(314), C(313), Z(314), C(314));
    I315 : HA port map (A(315), C(314), Z(315), C(315));
    I316 : HA port map (A(316), C(315), Z(316), C(316));
    I317 : HA port map (A(317), C(316), Z(317), C(317));
    I318 : HA port map (A(318), C(317), Z(318), C(318));
    I319 : HA port map (A(319), C(318), Z(319), C(319));
    I320 : HA port map (A(320), C(319), Z(320), C(320));
    I321 : HA port map (A(321), C(320), Z(321), C(321));
    I322 : HA port map (A(322), C(321), Z(322), C(322));
    I323 : HA port map (A(323), C(322), Z(323), C(323));
    I324 : HA port map (A(324), C(323), Z(324), C(324));
    I325 : HA port map (A(325), C(324), Z(325), C(325));
    I326 : HA port map (A(326), C(325), Z(326), C(326));
    I327 : HA port map (A(327), C(326), Z(327), C(327));
    I328 : HA port map (A(328), C(327), Z(328), C(328));
    I329 : HA port map (A(329), C(328), Z(329), C(329));
    I330 : HA port map (A(330), C(329), Z(330), C(330));
    I331 : HA port map (A(331), C(330), Z(331), C(331));
    I332 : HA port map (A(332), C(331), Z(332), C(332));
    I333 : HA port map (A(333), C(332), Z(333), C(333));
    I334 : HA port map (A(334), C(333), Z(334), C(334));
    I335 : HA port map (A(335), C(334), Z(335), C(335));
    I336 : HA port map (A(336), C(335), Z(336), C(336));
    I337 : HA port map (A(337), C(336), Z(337), C(337));
    I338 : HA port map (A(338), C(337), Z(338), C(338));
    I339 : HA port map (A(339), C(338), Z(339), C(339));
    I340 : HA port map (A(340), C(339), Z(340), C(340));
    I341 : HA port map (A(341), C(340), Z(341), C(341));
    I342 : HA port map (A(342), C(341), Z(342), C(342));
    I343 : HA port map (A(343), C(342), Z(343), C(343));
    I344 : HA port map (A(344), C(343), Z(344), C(344));
    I345 : HA port map (A(345), C(344), Z(345), C(345));
    I346 : HA port map (A(346), C(345), Z(346), C(346));
    I347 : HA port map (A(347), C(346), Z(347), C(347));
    I348 : HA port map (A(348), C(347), Z(348), C(348));
    I349 : HA port map (A(349), C(348), Z(349), C(349));
    I350 : HA port map (A(350), C(349), Z(350), C(350));
    I351 : HA port map (A(351), C(350), Z(351), C(351));
    I352 : HA port map (A(352), C(351), Z(352), C(352));
    I353 : HA port map (A(353), C(352), Z(353), C(353));
    I354 : HA port map (A(354), C(353), Z(354), C(354));
    I355 : HA port map (A(355), C(354), Z(355), C(355));
    I356 : HA port map (A(356), C(355), Z(356), C(356));
    I357 : HA port map (A(357), C(356), Z(357), C(357));
    I358 : HA port map (A(358), C(357), Z(358), C(358));
    I359 : HA port map (A(359), C(358), Z(359), C(359));
    I360 : HA port map (A(360), C(359), Z(360), C(360));
    I361 : HA port map (A(361), C(360), Z(361), C(361));
    I362 : HA port map (A(362), C(361), Z(362), C(362));
    I363 : HA port map (A(363), C(362), Z(363), C(363));
    I364 : HA port map (A(364), C(363), Z(364), C(364));
    I365 : HA port map (A(365), C(364), Z(365), C(365));
    I366 : HA port map (A(366), C(365), Z(366), C(366));
    I367 : HA port map (A(367), C(366), Z(367), C(367));
    I368 : HA port map (A(368), C(367), Z(368), C(368));
    I369 : HA port map (A(369), C(368), Z(369), C(369));
    I370 : HA port map (A(370), C(369), Z(370), C(370));
    I371 : HA port map (A(371), C(370), Z(371), C(371));
    I372 : HA port map (A(372), C(371), Z(372), C(372));
    I373 : HA port map (A(373), C(372), Z(373), C(373));
    I374 : HA port map (A(374), C(373), Z(374), C(374));
    I375 : HA port map (A(375), C(374), Z(375), C(375));
    I376 : HA port map (A(376), C(375), Z(376), C(376));
    I377 : HA port map (A(377), C(376), Z(377), C(377));
    I378 : HA port map (A(378), C(377), Z(378), C(378));
    I379 : HA port map (A(379), C(378), Z(379), C(379));
    I380 : HA port map (A(380), C(379), Z(380), C(380));
    I381 : HA port map (A(381), C(380), Z(381), C(381));
    I382 : HA port map (A(382), C(381), Z(382), C(382));
    I383 : HA port map (A(383), C(382), Z(383), C(383));
    I384 : HA port map (A(384), C(383), Z(384), C(384));
    I385 : HA port map (A(385), C(384), Z(385), C(385));
    I386 : HA port map (A(386), C(385), Z(386), C(386));
    I387 : HA port map (A(387), C(386), Z(387), C(387));
    I388 : HA port map (A(388), C(387), Z(388), C(388));
    I389 : HA port map (A(389), C(388), Z(389), C(389));
    I390 : HA port map (A(390), C(389), Z(390), C(390));
    I391 : HA port map (A(391), C(390), Z(391), C(391));
    I392 : HA port map (A(392), C(391), Z(392), C(392));
    I393 : HA port map (A(393), C(392), Z(393), C(393));
    I394 : HA port map (A(394), C(393), Z(394), C(394));
    I395 : HA port map (A(395), C(394), Z(395), C(395));
    I396 : HA port map (A(396), C(395), Z(396), C(396));
    I397 : HA port map (A(397), C(396), Z(397), C(397));
    I398 : HA port map (A(398), C(397), Z(398), C(398));
    I399 : HA port map (A(399), C(398), Z(399), C(399));
    I400 : HA port map (A(400), C(399), Z(400), C(400));
    I401 : HA port map (A(401), C(400), Z(401), C(401));
    I402 : HA port map (A(402), C(401), Z(402), C(402));
    I403 : HA port map (A(403), C(402), Z(403), C(403));
    I404 : HA port map (A(404), C(403), Z(404), C(404));
    I405 : HA port map (A(405), C(404), Z(405), C(405));
    I406 : HA port map (A(406), C(405), Z(406), C(406));
    I407 : HA port map (A(407), C(406), Z(407), C(407));
    I408 : HA port map (A(408), C(407), Z(408), C(408));
    I409 : HA port map (A(409), C(408), Z(409), C(409));
    I410 : HA port map (A(410), C(409), Z(410), C(410));
    I411 : HA port map (A(411), C(410), Z(411), C(411));
    I412 : HA port map (A(412), C(411), Z(412), C(412));
    I413 : HA port map (A(413), C(412), Z(413), C(413));
    I414 : HA port map (A(414), C(413), Z(414), C(414));
    I415 : HA port map (A(415), C(414), Z(415), C(415));
    I416 : HA port map (A(416), C(415), Z(416), C(416));
    I417 : HA port map (A(417), C(416), Z(417), C(417));
    I418 : HA port map (A(418), C(417), Z(418), C(418));
    I419 : HA port map (A(419), C(418), Z(419), C(419));
    I420 : HA port map (A(420), C(419), Z(420), C(420));
    I421 : HA port map (A(421), C(420), Z(421), C(421));
    I422 : HA port map (A(422), C(421), Z(422), C(422));
    I423 : HA port map (A(423), C(422), Z(423), C(423));
    I424 : HA port map (A(424), C(423), Z(424), C(424));
    I425 : HA port map (A(425), C(424), Z(425), C(425));
    I426 : HA port map (A(426), C(425), Z(426), C(426));
    I427 : HA port map (A(427), C(426), Z(427), C(427));
    I428 : HA port map (A(428), C(427), Z(428), C(428));
    I429 : HA port map (A(429), C(428), Z(429), C(429));
    I430 : HA port map (A(430), C(429), Z(430), C(430));
    I431 : HA port map (A(431), C(430), Z(431), C(431));
    I432 : HA port map (A(432), C(431), Z(432), C(432));
    I433 : HA port map (A(433), C(432), Z(433), C(433));
    I434 : HA port map (A(434), C(433), Z(434), C(434));
    I435 : HA port map (A(435), C(434), Z(435), C(435));
    I436 : HA port map (A(436), C(435), Z(436), C(436));
    I437 : HA port map (A(437), C(436), Z(437), C(437));
    I438 : HA port map (A(438), C(437), Z(438), C(438));
    I439 : HA port map (A(439), C(438), Z(439), C(439));
    I440 : HA port map (A(440), C(439), Z(440), C(440));
    I441 : HA port map (A(441), C(440), Z(441), C(441));
    I442 : HA port map (A(442), C(441), Z(442), C(442));
    I443 : HA port map (A(443), C(442), Z(443), C(443));
    I444 : HA port map (A(444), C(443), Z(444), C(444));
    I445 : HA port map (A(445), C(444), Z(445), C(445));
    I446 : HA port map (A(446), C(445), Z(446), C(446));
    I447 : HA port map (A(447), C(446), Z(447), C(447));
    I448 : HA port map (A(448), C(447), Z(448), C(448));
    I449 : HA port map (A(449), C(448), Z(449), C(449));
    I450 : HA port map (A(450), C(449), Z(450), C(450));
    I451 : HA port map (A(451), C(450), Z(451), C(451));
    I452 : HA port map (A(452), C(451), Z(452), C(452));
    I453 : HA port map (A(453), C(452), Z(453), C(453));
    I454 : HA port map (A(454), C(453), Z(454), C(454));
    I455 : HA port map (A(455), C(454), Z(455), C(455));
    I456 : HA port map (A(456), C(455), Z(456), C(456));
    I457 : HA port map (A(457), C(456), Z(457), C(457));
    I458 : HA port map (A(458), C(457), Z(458), C(458));
    I459 : HA port map (A(459), C(458), Z(459), C(459));
    I460 : HA port map (A(460), C(459), Z(460), C(460));
    I461 : HA port map (A(461), C(460), Z(461), C(461));
    I462 : HA port map (A(462), C(461), Z(462), C(462));
    I463 : HA port map (A(463), C(462), Z(463), C(463));
    I464 : HA port map (A(464), C(463), Z(464), C(464));
    I465 : HA port map (A(465), C(464), Z(465), C(465));
    I466 : HA port map (A(466), C(465), Z(466), C(466));
    I467 : HA port map (A(467), C(466), Z(467), C(467));
    I468 : HA port map (A(468), C(467), Z(468), C(468));
    I469 : HA port map (A(469), C(468), Z(469), C(469));
    I470 : HA port map (A(470), C(469), Z(470), C(470));
    I471 : HA port map (A(471), C(470), Z(471), C(471));
    I472 : HA port map (A(472), C(471), Z(472), C(472));
    I473 : HA port map (A(473), C(472), Z(473), C(473));
    I474 : HA port map (A(474), C(473), Z(474), C(474));
    I475 : HA port map (A(475), C(474), Z(475), C(475));
    I476 : HA port map (A(476), C(475), Z(476), C(476));
    I477 : HA port map (A(477), C(476), Z(477), C(477));
    I478 : HA port map (A(478), C(477), Z(478), C(478));
    I479 : HA port map (A(479), C(478), Z(479), C(479));
    I480 : HA port map (A(480), C(479), Z(480), C(480));
    I481 : HA port map (A(481), C(480), Z(481), C(481));
    I482 : HA port map (A(482), C(481), Z(482), C(482));
    I483 : HA port map (A(483), C(482), Z(483), C(483));
    I484 : HA port map (A(484), C(483), Z(484), C(484));
    I485 : HA port map (A(485), C(484), Z(485), C(485));
    I486 : HA port map (A(486), C(485), Z(486), C(486));
    I487 : HA port map (A(487), C(486), Z(487), C(487));
    I488 : HA port map (A(488), C(487), Z(488), C(488));
    I489 : HA port map (A(489), C(488), Z(489), C(489));
    I490 : HA port map (A(490), C(489), Z(490), C(490));
    I491 : HA port map (A(491), C(490), Z(491), C(491));
    I492 : HA port map (A(492), C(491), Z(492), C(492));
    I493 : HA port map (A(493), C(492), Z(493), C(493));
    I494 : HA port map (A(494), C(493), Z(494), C(494));
    I495 : HA port map (A(495), C(494), Z(495), C(495));
    I496 : HA port map (A(496), C(495), Z(496), C(496));
    I497 : HA port map (A(497), C(496), Z(497), C(497));
    I498 : HA port map (A(498), C(497), Z(498), C(498));
    I499 : HA port map (A(499), C(498), Z(499), C(499));
    I500 : HA port map (A(500), C(499), Z(500), C(500));
    I501 : HA port map (A(501), C(500), Z(501), C(501));
    I502 : HA port map (A(502), C(501), Z(502), C(502));
    I503 : HA port map (A(503), C(502), Z(503), C(503));
    I504 : HA port map (A(504), C(503), Z(504), C(504));
    I505 : HA port map (A(505), C(504), Z(505), C(505));
    I506 : HA port map (A(506), C(505), Z(506), C(506));
    I507 : HA port map (A(507), C(506), Z(507), C(507));
    I508 : HA port map (A(508), C(507), Z(508), C(508));
    I509 : HA port map (A(509), C(508), Z(509), C(509));
    I510 : HA port map (A(510), C(509), Z(510), C(510));
    I511 : HA port map (A(511), C(510), Z(511), C(511));
    I512 : HA port map (A(512), C(511), Z(512), C(512));
    I513 : HA port map (A(513), C(512), Z(513), C(513));
    I514 : HA port map (A(514), C(513), Z(514), C(514));
    I515 : HA port map (A(515), C(514), Z(515), C(515));
    I516 : HA port map (A(516), C(515), Z(516), C(516));
    I517 : HA port map (A(517), C(516), Z(517), C(517));
    I518 : HA port map (A(518), C(517), Z(518), C(518));
    I519 : HA port map (A(519), C(518), Z(519), C(519));
    I520 : HA port map (A(520), C(519), Z(520), C(520));
    I521 : HA port map (A(521), C(520), Z(521), C(521));
    I522 : HA port map (A(522), C(521), Z(522), C(522));
    I523 : HA port map (A(523), C(522), Z(523), C(523));
    I524 : HA port map (A(524), C(523), Z(524), C(524));
    I525 : HA port map (A(525), C(524), Z(525), C(525));
    I526 : HA port map (A(526), C(525), Z(526), C(526));
    I527 : HA port map (A(527), C(526), Z(527), C(527));
    I528 : HA port map (A(528), C(527), Z(528), C(528));
    I529 : HA port map (A(529), C(528), Z(529), C(529));
    I530 : HA port map (A(530), C(529), Z(530), C(530));
    I531 : HA port map (A(531), C(530), Z(531), C(531));
    I532 : HA port map (A(532), C(531), Z(532), C(532));
    I533 : HA port map (A(533), C(532), Z(533), C(533));
    I534 : HA port map (A(534), C(533), Z(534), C(534));
    I535 : HA port map (A(535), C(534), Z(535), C(535));
    I536 : HA port map (A(536), C(535), Z(536), C(536));
    I537 : HA port map (A(537), C(536), Z(537), C(537));
    I538 : HA port map (A(538), C(537), Z(538), C(538));
    I539 : HA port map (A(539), C(538), Z(539), C(539));
    I540 : HA port map (A(540), C(539), Z(540), C(540));
    I541 : HA port map (A(541), C(540), Z(541), C(541));
    I542 : HA port map (A(542), C(541), Z(542), C(542));
    I543 : HA port map (A(543), C(542), Z(543), C(543));
    I544 : HA port map (A(544), C(543), Z(544), C(544));
    I545 : HA port map (A(545), C(544), Z(545), C(545));
    I546 : HA port map (A(546), C(545), Z(546), C(546));
    I547 : HA port map (A(547), C(546), Z(547), C(547));
    I548 : HA port map (A(548), C(547), Z(548), C(548));
    I549 : HA port map (A(549), C(548), Z(549), C(549));
    I550 : HA port map (A(550), C(549), Z(550), C(550));
    I551 : HA port map (A(551), C(550), Z(551), C(551));
    I552 : HA port map (A(552), C(551), Z(552), C(552));
    I553 : HA port map (A(553), C(552), Z(553), C(553));
    I554 : HA port map (A(554), C(553), Z(554), C(554));
    I555 : HA port map (A(555), C(554), Z(555), C(555));
    I556 : HA port map (A(556), C(555), Z(556), C(556));
    I557 : HA port map (A(557), C(556), Z(557), C(557));
    I558 : HA port map (A(558), C(557), Z(558), C(558));
    I559 : HA port map (A(559), C(558), Z(559), C(559));
    I560 : HA port map (A(560), C(559), Z(560), C(560));
    I561 : HA port map (A(561), C(560), Z(561), C(561));
    I562 : HA port map (A(562), C(561), Z(562), C(562));
    I563 : HA port map (A(563), C(562), Z(563), C(563));
    I564 : HA port map (A(564), C(563), Z(564), C(564));
    I565 : HA port map (A(565), C(564), Z(565), C(565));
    I566 : HA port map (A(566), C(565), Z(566), C(566));
    I567 : HA port map (A(567), C(566), Z(567), C(567));
    I568 : HA port map (A(568), C(567), Z(568), C(568));
    I569 : HA port map (A(569), C(568), Z(569), C(569));
    I570 : HA port map (A(570), C(569), Z(570), C(570));
    I571 : HA port map (A(571), C(570), Z(571), C(571));
    I572 : HA port map (A(572), C(571), Z(572), C(572));
    I573 : HA port map (A(573), C(572), Z(573), C(573));
    I574 : HA port map (A(574), C(573), Z(574), C(574));
    I575 : HA port map (A(575), C(574), Z(575), C(575));
    I576 : HA port map (A(576), C(575), Z(576), C(576));
    I577 : HA port map (A(577), C(576), Z(577), C(577));
    I578 : HA port map (A(578), C(577), Z(578), C(578));
    I579 : HA port map (A(579), C(578), Z(579), C(579));
    I580 : HA port map (A(580), C(579), Z(580), C(580));
    I581 : HA port map (A(581), C(580), Z(581), C(581));
    I582 : HA port map (A(582), C(581), Z(582), C(582));
    I583 : HA port map (A(583), C(582), Z(583), C(583));
    I584 : HA port map (A(584), C(583), Z(584), C(584));
    I585 : HA port map (A(585), C(584), Z(585), C(585));
    I586 : HA port map (A(586), C(585), Z(586), C(586));
    I587 : HA port map (A(587), C(586), Z(587), C(587));
    I588 : HA port map (A(588), C(587), Z(588), C(588));
    I589 : HA port map (A(589), C(588), Z(589), C(589));
    I590 : HA port map (A(590), C(589), Z(590), C(590));
    I591 : HA port map (A(591), C(590), Z(591), C(591));
    I592 : HA port map (A(592), C(591), Z(592), C(592));
    I593 : HA port map (A(593), C(592), Z(593), C(593));
    I594 : HA port map (A(594), C(593), Z(594), C(594));
    I595 : HA port map (A(595), C(594), Z(595), C(595));
    I596 : HA port map (A(596), C(595), Z(596), C(596));
    I597 : HA port map (A(597), C(596), Z(597), C(597));
    I598 : HA port map (A(598), C(597), Z(598), C(598));
    I599 : HA port map (A(599), C(598), Z(599), C(599));
    I600 : HA port map (A(600), C(599), Z(600), C(600));
    I601 : HA port map (A(601), C(600), Z(601), C(601));
    I602 : HA port map (A(602), C(601), Z(602), C(602));
    I603 : HA port map (A(603), C(602), Z(603), C(603));
    I604 : HA port map (A(604), C(603), Z(604), C(604));
    I605 : HA port map (A(605), C(604), Z(605), C(605));
    I606 : HA port map (A(606), C(605), Z(606), C(606));
    I607 : HA port map (A(607), C(606), Z(607), C(607));
    I608 : HA port map (A(608), C(607), Z(608), C(608));
    I609 : HA port map (A(609), C(608), Z(609), C(609));
    I610 : HA port map (A(610), C(609), Z(610), C(610));
    I611 : HA port map (A(611), C(610), Z(611), C(611));
    I612 : HA port map (A(612), C(611), Z(612), C(612));
    I613 : HA port map (A(613), C(612), Z(613), C(613));
    I614 : HA port map (A(614), C(613), Z(614), C(614));
    I615 : HA port map (A(615), C(614), Z(615), C(615));
    I616 : HA port map (A(616), C(615), Z(616), C(616));
    I617 : HA port map (A(617), C(616), Z(617), C(617));
    I618 : HA port map (A(618), C(617), Z(618), C(618));
    I619 : HA port map (A(619), C(618), Z(619), C(619));
    I620 : HA port map (A(620), C(619), Z(620), C(620));
    I621 : HA port map (A(621), C(620), Z(621), C(621));
    I622 : HA port map (A(622), C(621), Z(622), C(622));
    I623 : HA port map (A(623), C(622), Z(623), C(623));
    I624 : HA port map (A(624), C(623), Z(624), C(624));
    I625 : HA port map (A(625), C(624), Z(625), C(625));
    I626 : HA port map (A(626), C(625), Z(626), C(626));
    I627 : HA port map (A(627), C(626), Z(627), C(627));
    I628 : HA port map (A(628), C(627), Z(628), C(628));
    I629 : HA port map (A(629), C(628), Z(629), C(629));
    I630 : HA port map (A(630), C(629), Z(630), C(630));
    I631 : HA port map (A(631), C(630), Z(631), C(631));
    I632 : HA port map (A(632), C(631), Z(632), C(632));
    I633 : HA port map (A(633), C(632), Z(633), C(633));
    I634 : HA port map (A(634), C(633), Z(634), C(634));
    I635 : HA port map (A(635), C(634), Z(635), C(635));
    I636 : HA port map (A(636), C(635), Z(636), C(636));
    I637 : HA port map (A(637), C(636), Z(637), C(637));
    I638 : HA port map (A(638), C(637), Z(638), C(638));
    I639 : HA port map (A(639), C(638), Z(639), C(639));
    I640 : HA port map (A(640), C(639), Z(640), C(640));
    I641 : HA port map (A(641), C(640), Z(641), C(641));
    I642 : HA port map (A(642), C(641), Z(642), C(642));
    I643 : HA port map (A(643), C(642), Z(643), C(643));
    I644 : HA port map (A(644), C(643), Z(644), C(644));
    I645 : HA port map (A(645), C(644), Z(645), C(645));
    I646 : HA port map (A(646), C(645), Z(646), C(646));
    I647 : HA port map (A(647), C(646), Z(647), C(647));
    I648 : HA port map (A(648), C(647), Z(648), C(648));
    I649 : HA port map (A(649), C(648), Z(649), C(649));
    I650 : HA port map (A(650), C(649), Z(650), C(650));
    I651 : HA port map (A(651), C(650), Z(651), C(651));
    I652 : HA port map (A(652), C(651), Z(652), C(652));
    I653 : HA port map (A(653), C(652), Z(653), C(653));
    I654 : HA port map (A(654), C(653), Z(654), C(654));
    I655 : HA port map (A(655), C(654), Z(655), C(655));
    I656 : HA port map (A(656), C(655), Z(656), C(656));
    I657 : HA port map (A(657), C(656), Z(657), C(657));
    I658 : HA port map (A(658), C(657), Z(658), C(658));
    I659 : HA port map (A(659), C(658), Z(659), C(659));
    I660 : HA port map (A(660), C(659), Z(660), C(660));
    I661 : HA port map (A(661), C(660), Z(661), C(661));
    I662 : HA port map (A(662), C(661), Z(662), C(662));
    I663 : HA port map (A(663), C(662), Z(663), C(663));
    I664 : HA port map (A(664), C(663), Z(664), C(664));
    I665 : HA port map (A(665), C(664), Z(665), C(665));
    I666 : HA port map (A(666), C(665), Z(666), C(666));
    I667 : HA port map (A(667), C(666), Z(667), C(667));
    I668 : HA port map (A(668), C(667), Z(668), C(668));
    I669 : HA port map (A(669), C(668), Z(669), C(669));
    I670 : HA port map (A(670), C(669), Z(670), C(670));
    I671 : HA port map (A(671), C(670), Z(671), C(671));
    I672 : HA port map (A(672), C(671), Z(672), C(672));
    I673 : HA port map (A(673), C(672), Z(673), C(673));
    I674 : HA port map (A(674), C(673), Z(674), C(674));
    I675 : HA port map (A(675), C(674), Z(675), C(675));
    I676 : HA port map (A(676), C(675), Z(676), C(676));
    I677 : HA port map (A(677), C(676), Z(677), C(677));
    I678 : HA port map (A(678), C(677), Z(678), C(678));
    I679 : HA port map (A(679), C(678), Z(679), C(679));
    I680 : HA port map (A(680), C(679), Z(680), C(680));
    I681 : HA port map (A(681), C(680), Z(681), C(681));
    I682 : HA port map (A(682), C(681), Z(682), C(682));
    I683 : HA port map (A(683), C(682), Z(683), C(683));
    I684 : HA port map (A(684), C(683), Z(684), C(684));
    I685 : HA port map (A(685), C(684), Z(685), C(685));
    I686 : HA port map (A(686), C(685), Z(686), C(686));
    I687 : HA port map (A(687), C(686), Z(687), C(687));
    I688 : HA port map (A(688), C(687), Z(688), C(688));
    I689 : HA port map (A(689), C(688), Z(689), C(689));
    I690 : HA port map (A(690), C(689), Z(690), C(690));
    I691 : HA port map (A(691), C(690), Z(691), C(691));
    I692 : HA port map (A(692), C(691), Z(692), C(692));
    I693 : HA port map (A(693), C(692), Z(693), C(693));
    I694 : HA port map (A(694), C(693), Z(694), C(694));
    I695 : HA port map (A(695), C(694), Z(695), C(695));
    I696 : HA port map (A(696), C(695), Z(696), C(696));
    I697 : HA port map (A(697), C(696), Z(697), C(697));
    I698 : HA port map (A(698), C(697), Z(698), C(698));
    I699 : HA port map (A(699), C(698), Z(699), C(699));
    I700 : HA port map (A(700), C(699), Z(700), C(700));
    I701 : HA port map (A(701), C(700), Z(701), C(701));
    I702 : HA port map (A(702), C(701), Z(702), C(702));
    I703 : HA port map (A(703), C(702), Z(703), C(703));
    I704 : HA port map (A(704), C(703), Z(704), C(704));
    I705 : HA port map (A(705), C(704), Z(705), C(705));
    I706 : HA port map (A(706), C(705), Z(706), C(706));
    I707 : HA port map (A(707), C(706), Z(707), C(707));
    I708 : HA port map (A(708), C(707), Z(708), C(708));
    I709 : HA port map (A(709), C(708), Z(709), C(709));
    I710 : HA port map (A(710), C(709), Z(710), C(710));
    I711 : HA port map (A(711), C(710), Z(711), C(711));
    I712 : HA port map (A(712), C(711), Z(712), C(712));
    I713 : HA port map (A(713), C(712), Z(713), C(713));
    I714 : HA port map (A(714), C(713), Z(714), C(714));
    I715 : HA port map (A(715), C(714), Z(715), C(715));
    I716 : HA port map (A(716), C(715), Z(716), C(716));
    I717 : HA port map (A(717), C(716), Z(717), C(717));
    I718 : HA port map (A(718), C(717), Z(718), C(718));
    I719 : HA port map (A(719), C(718), Z(719), C(719));
    I720 : HA port map (A(720), C(719), Z(720), C(720));
    I721 : HA port map (A(721), C(720), Z(721), C(721));
    I722 : HA port map (A(722), C(721), Z(722), C(722));
    I723 : HA port map (A(723), C(722), Z(723), C(723));
    I724 : HA port map (A(724), C(723), Z(724), C(724));
    I725 : HA port map (A(725), C(724), Z(725), C(725));
    I726 : HA port map (A(726), C(725), Z(726), C(726));
    I727 : HA port map (A(727), C(726), Z(727), C(727));
    I728 : HA port map (A(728), C(727), Z(728), C(728));
    I729 : HA port map (A(729), C(728), Z(729), C(729));
    I730 : HA port map (A(730), C(729), Z(730), C(730));
    I731 : HA port map (A(731), C(730), Z(731), C(731));
    I732 : HA port map (A(732), C(731), Z(732), C(732));
    I733 : HA port map (A(733), C(732), Z(733), C(733));
    I734 : HA port map (A(734), C(733), Z(734), C(734));
    I735 : HA port map (A(735), C(734), Z(735), C(735));
    I736 : HA port map (A(736), C(735), Z(736), C(736));
    I737 : HA port map (A(737), C(736), Z(737), C(737));
    I738 : HA port map (A(738), C(737), Z(738), C(738));
    I739 : HA port map (A(739), C(738), Z(739), C(739));
    I740 : HA port map (A(740), C(739), Z(740), C(740));
    I741 : HA port map (A(741), C(740), Z(741), C(741));
    I742 : HA port map (A(742), C(741), Z(742), C(742));
    I743 : HA port map (A(743), C(742), Z(743), C(743));
    I744 : HA port map (A(744), C(743), Z(744), C(744));
    I745 : HA port map (A(745), C(744), Z(745), C(745));
    I746 : HA port map (A(746), C(745), Z(746), C(746));
    I747 : HA port map (A(747), C(746), Z(747), C(747));
    I748 : HA port map (A(748), C(747), Z(748), C(748));
    I749 : HA port map (A(749), C(748), Z(749), C(749));
    I750 : HA port map (A(750), C(749), Z(750), C(750));
    I751 : HA port map (A(751), C(750), Z(751), C(751));
    I752 : HA port map (A(752), C(751), Z(752), C(752));
    I753 : HA port map (A(753), C(752), Z(753), C(753));
    I754 : HA port map (A(754), C(753), Z(754), C(754));
    I755 : HA port map (A(755), C(754), Z(755), C(755));
    I756 : HA port map (A(756), C(755), Z(756), C(756));
    I757 : HA port map (A(757), C(756), Z(757), C(757));
    I758 : HA port map (A(758), C(757), Z(758), C(758));
    I759 : HA port map (A(759), C(758), Z(759), C(759));
    I760 : HA port map (A(760), C(759), Z(760), C(760));
    I761 : HA port map (A(761), C(760), Z(761), C(761));
    I762 : HA port map (A(762), C(761), Z(762), C(762));
    I763 : HA port map (A(763), C(762), Z(763), C(763));
    I764 : HA port map (A(764), C(763), Z(764), C(764));
    I765 : HA port map (A(765), C(764), Z(765), C(765));
    I766 : HA port map (A(766), C(765), Z(766), C(766));
    I767 : HA port map (A(767), C(766), Z(767), C(767));
    I768 : HA port map (A(768), C(767), Z(768), C(768));
    I769 : HA port map (A(769), C(768), Z(769), C(769));
    I770 : HA port map (A(770), C(769), Z(770), C(770));
    I771 : HA port map (A(771), C(770), Z(771), C(771));
    I772 : HA port map (A(772), C(771), Z(772), C(772));
    I773 : HA port map (A(773), C(772), Z(773), C(773));
    I774 : HA port map (A(774), C(773), Z(774), C(774));
    I775 : HA port map (A(775), C(774), Z(775), C(775));
    I776 : HA port map (A(776), C(775), Z(776), C(776));
    I777 : HA port map (A(777), C(776), Z(777), C(777));
    I778 : HA port map (A(778), C(777), Z(778), C(778));
    I779 : HA port map (A(779), C(778), Z(779), C(779));
    I780 : HA port map (A(780), C(779), Z(780), C(780));
    I781 : HA port map (A(781), C(780), Z(781), C(781));
    I782 : HA port map (A(782), C(781), Z(782), C(782));
    I783 : HA port map (A(783), C(782), Z(783), C(783));
    I784 : HA port map (A(784), C(783), Z(784), C(784));
    I785 : HA port map (A(785), C(784), Z(785), C(785));
    I786 : HA port map (A(786), C(785), Z(786), C(786));
    I787 : HA port map (A(787), C(786), Z(787), C(787));
    I788 : HA port map (A(788), C(787), Z(788), C(788));
    I789 : HA port map (A(789), C(788), Z(789), C(789));
    I790 : HA port map (A(790), C(789), Z(790), C(790));
    I791 : HA port map (A(791), C(790), Z(791), C(791));
    I792 : HA port map (A(792), C(791), Z(792), C(792));
    I793 : HA port map (A(793), C(792), Z(793), C(793));
    I794 : HA port map (A(794), C(793), Z(794), C(794));
    I795 : HA port map (A(795), C(794), Z(795), C(795));
    I796 : HA port map (A(796), C(795), Z(796), C(796));
    I797 : HA port map (A(797), C(796), Z(797), C(797));
    I798 : HA port map (A(798), C(797), Z(798), C(798));
    I799 : HA port map (A(799), C(798), Z(799), C(799));
 

	 
END ARC;

